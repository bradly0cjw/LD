module tb_Decoder(
    reg A
)
endmodule
